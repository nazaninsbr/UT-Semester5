library verilog;
use verilog.vl_types.all;
entity test_Seg is
end test_Seg;
