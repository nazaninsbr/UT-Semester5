library verilog;
use verilog.vl_types.all;
entity test_clockDivider is
end test_clockDivider;
