library verilog;
use verilog.vl_types.all;
entity test_pwm is
end test_pwm;
