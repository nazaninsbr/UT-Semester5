module part1(); 

endmodule 