library verilog;
use verilog.vl_types.all;
entity test_comparator is
end test_comparator;
